class mem_common;

  static int num_matches;
  static int num_mismatches;
endclass
